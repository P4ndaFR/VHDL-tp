---___      ___ ___  ___  ________  ___
--|\  \    /  /|\  \|\  \|\   ___ \|\  \
--\ \  \  /  / | \  \\\  \ \  \_|\ \ \  \
-- \ \  \/  / / \ \   __  \ \  \ \\ \ \  \
--  \ \    / /   \ \  \ \  \ \  \_\\ \ \  \____
--   \ \__/ /     \ \__\ \__\ \_______\ \_______\
--    \|__|/       \|__|\|__|\|_______|\|_______|
-------------------------------------------------
-- Fichier comparateur.vhd
-- Antoine Blondeau
-- comparaison de 2 nombres sur 4 bits
-------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity trans_hexa_7seg is
  port
  (
    code_e: in std_logic_vector( 3 downto 0 );
    code_s: out std_logic_vector( 6 downto 0 )
  );
end trans_hexa_7seg;
architecture beh of trans_hexa_7seg is
  begin
    with code_e select
    code_s <=
    "1000000" when "0000",  --0
    "1111001" when "0001",  --1
    "0100100" when "0010",  --2
    "0110000" when "0011",  --3
    "0011001" when "0100",  --4
    "0010010" when "0101",  --5
    "0000010" when "0110",  --6
    "1111000" when "0111",  --7
    "0000000" when "1000",  --8
    "0010000" when "1001",  --9
    "1111111" when others;  --else
end beh;
